package common_constants;
    parameter AXI_BURST_TYPE_INCR = 2'b01;
    parameter VGA_VISIBLE_WIDTH = 640;
    parameter VGA_VISIBLE_HEIGHT = 480;
    parameter DISP_ADDR_WIDTH = 30;
endpackage
